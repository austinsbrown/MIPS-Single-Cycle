`include "program_counter.v"
`include "instruction_memory.v"
`include "control.v"
`include "registers.v"

module datapath
(
    
);

    

endmodule